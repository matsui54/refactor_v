module foo(
  AAA,
  BBB,
  CCC,
  DDD,
  EEE
);
  input AAA;
  input BBB;
  input CCC;
  input DDD;
  output EEE;
endmodule
