// ======================================================
// bar.sv : 1行1宣言のポート宣言（出力がベクタ）
// ======================================================
module bar(
  P,
  Q,
  R,
  S
);
  input  [15:0] P;
  input         Q;
  output [15:0] R;
  output [7:0]  S;

  // テスト用の簡単な出力計算
  assign R = Q ? {P[7:0], P[15:8]} : P;
  assign S = P[7:0] ^ P[15:8];
endmodule
